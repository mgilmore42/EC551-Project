`ifndef _my_incl_vh_
    `define _my_incl_vh_
    `define dwidth_dat 12
    `define dwidth_slice 5
    `define dwss 25 // must be dwidth_slice**2
    `define dwidth_kernel 8
    `define dwidth_div 4
    `define awidth_pbuff 10
    `define awidth_fbuff 19
    `define hwidth 640
    `define vwidth 480
`endif
