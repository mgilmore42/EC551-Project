`ifndef _my_incl_vh_
    `define _my_incl_vh_
    `define dwidth_dat 12
    `define dwidth_slice 9
    `define awidth_pbuff 10
    `define awidth_fbuff 19
    `define hwidth 640
    `define vwidth 480
//    `define dwidth_dat 16
//    `define awidth_mem 12
//    `define awidth_reg 6
//    `define inst_start 31
//    `define clk_div 10
`endif
